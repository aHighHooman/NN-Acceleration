module matrixMultiplierSmall (
    input  logic        clk,
    input  logic        rst_n,
    input  logic signed [15:0] matrixA [3][3],
    input  logic signed [15:0] matrixB [3][3],
    output logic signed [31:0] resultMatrix [3][3]
);
    
endmodule